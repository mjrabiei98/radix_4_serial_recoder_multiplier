library verilog;
use verilog.vl_types.all;
entity recoder is
    port(
        x_1             : in     vl_logic;
        x_0             : in     vl_logic;
        c_in            : in     vl_logic;
        one             : in     vl_logic;
        neg             : in     vl_logic;
        zero            : in     vl_logic;
        c_out           : in     vl_logic
    );
end recoder;
